module wallData (   input [9:0]	addr,
					output [415:0]	data
				);

    parameter SIZE =  416;
    parameter BYTES_NO = 10;

    //wall sprite
	parameter [0:2**BYTES_NO-1][SIZE-1:0] WallSprite = {
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001111111111111111111111111111110010000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111110010000000000000000000000000000000000000000000000000000000000001001111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000001001111111111111111111111111111110010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000111100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000111100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001111111111111111111111111111110010000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111110010000000000000000000000000000000000000000000000000000000000001001111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000001001111111111111111111111111111110010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110010000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000001001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110010000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000010011111111111111111111111111111111111111111111111111111111111111001000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001111000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000011110000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010011111111111111111111111111111111111111111111111111111111111111001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000,


416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
416'b 00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001111111111111111111111111111110010000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111110010000000000000000000000000000000000000000000000000000000000001001111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000001001111111111111111111111111111110010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000111100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000111100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001001111111111111111111111111111110010000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111110010000000000000000000000000000000000000000000000000000000000001001111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000001001111111111111111111111111111110010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110010000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000001001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110010000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000010011111111111111111111111111111111111111111111111111111111111111001000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001111000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000011110000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010011111111111111111111111111111111111111111111111111111111111111001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000100111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000,
416'b 00000000000000100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000,
416'b 00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000


};

	assign data = WallSprite[addr];

endmodule 